-- Elementos de Sistemas
-- by Luciano Soares
-- HalfAdder.vhd

-- Implementa Half Adder

Library ieee;
use ieee.std_logic_1164.all;

entity HalfAdder is
	port(
		a,b:         in STD_LOGIC;   -- entradas
		soma,vaium: out STD_LOGIC   -- sum e carry
	);
end entity;

architecture rtl of HalfAdder is
  -- Aqui declaramos sinais (fios auxiliares)
  -- e componentes (outros módulos) que serao
  -- utilizados nesse modulo.


begin
  -- Implementação vem aqui!
  --u1: HalfAdder port map(a => SW(0), b => SW(1), soma => LEDR(0), vaium => LEDR(1));
  soma <= a xor b;
  vaium <= a and b;


end rtl;
